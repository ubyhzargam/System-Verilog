// Simple code to print all the elements of an array 

module tb;
  bit arr[]={1,0,1,1,1};
  initial
    begin
      $display("%p",arr);
    end
endmodule
